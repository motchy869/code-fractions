package main_pkg;
    parameter int BIT_WIDTH_REG_1 = 3;
    parameter int BIT_WIDTH_REG_2 = 8;
endpackage
