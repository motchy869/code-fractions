`ifdef MACROS_SVH_INCLUDED

`undef INCR_NON_BLK

`endif
