`ifndef MACROS_SVH_INCLUDED
`define MACROS_SVH_INCLUDED

`define INCR_NON_BLK(x,d=1) x <= x + $bits(x)'(d);

`endif
