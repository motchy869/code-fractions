package main_pkg;
    parameter BIT_WIDTH_REG_1 = 3;
    parameter BIT_WIDTH_REG_2 = 8;
endpackage
